/* Copyright(C) 2020 Cobac.Net All Rights Reserved. */
/* chapter: ��9�͉ۑ�       */
/* project: display_xga     */
/* outline: XGA�p�p�����[�^ */

/* XGA(1024�~768)�p�����[�^ */
localparam HPERIOD = 11'd1344;
localparam HFRONT  = 11'd24;
localparam HWIDTH  = 11'd136;
localparam HBACK   = 11'd160;

localparam VPERIOD = 10'd806;
localparam VFRONT  = 10'd3;
localparam VWIDTH  = 10'd6;
localparam VBACK   = 10'd29;
